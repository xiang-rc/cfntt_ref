module tf_ROM 
    #(parameter addr_rom_width = 9,
                 data_width = 42,
                 depth_rom = 341)
    (
    input clk,
    input [addr_rom_width-1:0] A,
    input REN,
    output reg [data_width-1:0] Q);
    
    always@(posedge clk)
    begin
    if(REN == 1'b1) begin
    case(A)
    9'd0: Q <= 42'b011011111001111010100011101000111111001011;
    9'd1: Q <= 42'b001101110101101010101110100010100110010011;
    9'd2: Q <= 42'b101001100100110101100110100010001001010001;
    9'd3: Q <= 42'b100110000100000000101101001001011011100100;
    9'd4: Q <= 42'b001100011110110111111101101100100111110001;
    9'd5: Q <= 42'b001001000011110111010010110000110000010011;
    9'd6: Q <= 42'b100011100000001001011100000010010000010110;
    9'd7: Q <= 42'b101100010001100010100100111110110000011001;
    9'd8: Q <= 42'b010011110111101011000100110000101110010011;
    9'd9: Q <= 42'b001100000100110101100110000010001110000000;
    9'd10: Q <= 42'b100100011011100100111001111110101101101111;
    9'd11: Q <= 42'b011111001000010111100001001010101011010011;
    9'd12: Q <= 42'b100100000101100101101100010000001110111011;
    9'd13: Q <= 42'b010010111011101011011100111010111101110101;
    9'd14: Q <= 42'b010010110001011001000100001101111101100010;
    9'd15: Q <= 42'b100011110000101001000110001010110100101011;
    9'd16: Q <= 42'b101011110110111001010100100100011001100011;
    9'd17: Q <= 42'b101011011010001000110000000110001111000010;
    9'd18: Q <= 42'b101111011101010111001000111110001000100000;
    9'd19: Q <= 42'b101001100111100110010111000001110100010011;
    9'd20: Q <= 42'b011101111111100001010100011100010000100110;
    9'd21: Q <= 42'b001001011000010001001110110000100001110110;
    9'd22: Q <= 42'b000001100001100100100001100010111111111110;
    9'd23: Q <= 42'b011100000101000100010010010001110011001010;
    9'd24: Q <= 42'b100001000010000110011000011000000010100000;
    9'd25: Q <= 42'b000011111110010001111101110101110001001111;
    9'd26: Q <= 42'b000000000110110000101101100101110011100010;
    9'd27: Q <= 42'b000110011000001000110010100000101001010101;
    9'd28: Q <= 42'b100001010011100011001010100101101110110110;
    9'd29: Q <= 42'b000001011000100010010111101010101001101111;
    9'd30: Q <= 42'b010011100101000001011001010001001101001010;
    9'd31: Q <= 42'b100100101000010000010100111010100100010000;
    9'd32: Q <= 42'b001011001010110001101010000001101101010110;
    9'd33: Q <= 42'b000110000000010010110100000100111111011001;
    9'd34: Q <= 42'b100101100010110111000001110101111011000011;
    9'd35: Q <= 42'b010010011010100011001101010010001011011101;
    9'd36: Q <= 42'b010011100110111001111101100010011110000011;
    9'd37: Q <= 42'b001000011101101001001110011100001111111001;
    9'd38: Q <= 42'b101111011000010000111111111010000101001110;
    9'd39: Q <= 42'b101111100100000000011110000001110000100101;
    9'd40: Q <= 42'b101111111111100000000000100110111111100110;
    9'd41: Q <= 42'b001101001001001010010111100000000110000110;
    9'd42: Q <= 42'b100100111000100110110010111000000110111010;
    9'd43: Q <= 42'b001111110110010100001011011000111011000010;
    9'd44: Q <= 42'b001000011111100111001000010001001111101101;
    9'd45: Q <= 42'b001110001101001001100101110110010110001011;
    9'd46: Q <= 42'b101010011011110101101001111100000011110010;
    9'd47: Q <= 42'b010100101010110000010101001110110111100000;
    9'd48: Q <= 42'b000110011111110000100010000001110110010111;
    9'd49: Q <= 42'b011100010011110111111011000010010010100001;
    9'd50: Q <= 42'b010100010010110001010110010110011001010000;
    9'd51: Q <= 42'b001111110101011000100000000110111010011111;
    9'd52: Q <= 42'b011100111000101001100010010010010011010110;
    9'd53: Q <= 42'b000011111010101000011001001110011010100010;
    9'd54: Q <= 42'b011100100100011010010010001000101111001000;
    9'd55: Q <= 42'b010011111000000110111100011010001111000001;
    9'd56: Q <= 42'b100001001111011000011000011000101110111000;
    9'd57: Q <= 42'b101011110110000011100011010110011010111111;
    9'd58: Q <= 42'b000100100100000000001001000110010110000011;
    9'd59: Q <= 42'b101110011011010011011000001100110110110110;
    9'd60: Q <= 42'b101011010010100110100101101100111110001010;
    9'd61: Q <= 42'b100110011111000011010011011000111110010001;
    9'd62: Q <= 42'b100101111110111001100000110100000110100100;
    9'd63: Q <= 42'b010111100001101011101001111000000111011100;
    9'd64: Q <= 42'b011000011010100111110111101000100010000010;
    9'd65: Q <= 42'b000001111011011001010101011001010100011111;
    9'd66: Q <= 42'b011111000100000111001110011110010010111101;
    9'd67: Q <= 42'b011010101111011000001010010110100110100011;
    9'd68: Q <= 42'b000101011000100110001110101000100011001001;
    9'd69: Q <= 42'b100011010100101011000100100010011001111100;
    9'd70: Q <= 42'b100110101111110000110011101101100001101010;
    9'd71: Q <= 42'b100000011101111000010101110100101110101011;
    9'd72: Q <= 42'b010100110101000101101000011100101000000110;
    9'd73: Q <= 42'b100110101000100011110110110100010010010000;
    9'd74: Q <= 42'b100100010010010100010110010000100001011111;
    9'd75: Q <= 42'b011011101110101000110010000100110010110000;
    9'd76: Q <= 42'b001011110010000010010101110000000110010100;
    9'd77: Q <= 42'b000110010111100010011010110001001111100000;
    9'd78: Q <= 42'b101011100000000010001001010110100110111010;
    9'd79: Q <= 42'b010101000111110000000111011010110000010111;
    9'd80: Q <= 42'b100111001110000111000011011000111011000100;
    9'd81: Q <= 42'b011010010010100111101111111101101010111101;
    9'd82: Q <= 42'b001111100100010010110001010110111001001110;
    9'd83: Q <= 42'b100111011111110000001000001010111000010100;
    9'd84: Q <= 42'b001101110010110110110000001110101010011111;
    9'd85: Q <= 42'b000000000001110000000011000100000101010111;
    9'd86: Q <= 42'b001100010100100101110001101100010010111000;
    9'd87: Q <= 42'b000011010011010001001110111110100010001101;
    9'd88: Q <= 42'b001100110101010001011100101101010001011011;
    9'd89: Q <= 42'b001100001100000001011110100010101000000001;
    9'd90: Q <= 42'b100000100111001010001110101000001011001101;
    9'd91: Q <= 42'b011000001110110000010101111001111111111010;
    9'd92: Q <= 42'b001101110100000101010000011110101010100100;
    9'd93: Q <= 42'b000000110110001001100011110100001011001100;
    9'd94: Q <= 42'b000010111111111010011101001000100110010010;
    9'd95: Q <= 42'b011010011010111010100011000001101011011001;
    9'd96: Q <= 42'b100111010111000110001100101100000110100000;
    9'd97: Q <= 42'b001100100111010101001111100110001100110011;
    9'd98: Q <= 42'b000101000000101000110111111110111001001011;
    9'd99: Q <= 42'b101001010101111001111111100001101011011101;
    9'd100: Q <= 42'b000111111001010100011000110110101100111111;
    9'd101: Q <= 42'b100010011101000010111101011010000001111010;
    9'd102: Q <= 42'b010010010101010010010011100101111001101000;
    9'd103: Q <= 42'b011110101001100100000001001100110000001111;
    9'd104: Q <= 42'b100111000011001010001100111010101001111000;
    9'd105: Q <= 42'b101011000000010011110111101100101010011101;
    9'd106: Q <= 42'b101100011110010101111111111000100011010100;
    9'd107: Q <= 42'b101111111010010000100100000010101000000010;
    9'd108: Q <= 42'b011010010101101001100111001001100100110101;
    9'd109: Q <= 42'b000111000010100010110101110001001111101110;
    9'd110: Q <= 42'b011110110001100011010110101001001101100011;
    9'd111: Q <= 42'b010011111011110000001101101001100100101100;
    9'd112: Q <= 42'b000100110001111000100011100010011000100001;
    9'd113: Q <= 42'b000011011100010001111010001000001111110110;
    9'd114: Q <= 42'b010101010101011001001011111100111000010111;
    9'd115: Q <= 42'b000011111101111001111111111001110011000101;
    9'd116: Q <= 42'b001010010011011010001111010010000010011011;
    9'd117: Q <= 42'b001111011010001001010100111100110100011111;
    9'd118: Q <= 42'b001000011110110110011001101010100001111001;
    9'd119: Q <= 42'b010101111001000110010001010100010001000100;
    9'd120: Q <= 42'b101011000100000010100101111110000110100011;
    9'd121: Q <= 42'b100100100001001010000100101001111110000011;
    9'd122: Q <= 42'b001110111111010000010101101101000010000011;
    9'd123: Q <= 42'b011001111000111000010101010010111110000100;
    9'd124: Q <= 42'b001100100101010010110110110101111101110011;
    9'd125: Q <= 42'b100100100000001001000100000000010001110000;
    9'd126: Q <= 42'b100011011000010000001010111000101101101110;
    9'd127: Q <= 42'b001010010010010001101001110110001101011011;
    9'd128: Q <= 42'b010010111101110000101101001101111001111000;
    9'd129: Q <= 42'b001111110100101000110000111001011111101111;
    9'd130: Q <= 42'b101100001011010001110100001010011111101101;
    9'd131: Q <= 42'b000011010011001011100101011110001110100110;
    9'd132: Q <= 42'b010001111011100100101001001001111011001101;
    9'd133: Q <= 42'b010010010011000011111001011100100011100011;
    9'd134: Q <= 42'b011100100001101001010011001010101000010011;
    9'd135: Q <= 42'b011011111100101000001000000001011000010101;
    9'd136: Q <= 42'b001110010101100000001001110001110000111010;
    9'd137: Q <= 42'b010101111100100011101011110001001011111100;
    9'd138: Q <= 42'b010011101100110101110001010001010110000100;
    9'd139: Q <= 42'b010110100111010000011010001010101110010110;
    9'd140: Q <= 42'b001100000100101011100011110000010010011000;
    9'd141: Q <= 42'b000010010000100010001110100100110110100111;
    9'd142: Q <= 42'b011101110011001010000001001000111101111001;
    9'd143: Q <= 42'b101110001111110101101111010010011111110000;
    9'd144: Q <= 42'b100101110000110101001101010100011011011100;
    9'd145: Q <= 42'b001011111110010101010011010100001001000011;
    9'd146: Q <= 42'b011000111101010111011000000000110000101010;
    9'd147: Q <= 42'b011001101110100111010101101101011101100011;
    9'd148: Q <= 42'b011101100100100001010000110101011101001110;
    9'd149: Q <= 42'b000001010101110110111000100010001001110100;
    9'd150: Q <= 42'b011011101001100111111011100010011100001100;
    9'd151: Q <= 42'b010001101110101001001001100110001010100111;
    9'd152: Q <= 42'b000100101110001000111100101001110110101100;
    9'd153: Q <= 42'b010101001001000100111100000100001101110001;
    9'd154: Q <= 42'b001101101110110100101010110000101001001101;
    9'd155: Q <= 42'b100011001100110100100101101010100001111010;
    9'd156: Q <= 42'b000100110000101000101000110001101010101100;
    9'd157: Q <= 42'b101001010110000110101010010101111011000110;
    9'd158: Q <= 42'b000010110011001000100110011100011000010011;
    9'd159: Q <= 42'b101110011000010000111111001010011011100011;
    9'd160: Q <= 42'b001000011101000000110001001101110000010010;
    9'd161: Q <= 42'b101010000000011011110100000110111111101001;
    9'd162: Q <= 42'b000101010111010100110011000010011001001100;
    9'd163: Q <= 42'b001001011111010001010010100100010100000000;
    9'd164: Q <= 42'b000010110011011010000000000001010110101011;
    9'd165: Q <= 42'b001000000100011011111100011100110000110000;
    9'd166: Q <= 42'b100010001100110011011100110000110111010000;
    9'd167: Q <= 42'b001101101001111011110001000001011000001110;
    9'd168: Q <= 42'b101001001001011011000001011000111101100101;
    9'd169: Q <= 42'b101011000001100011011001010100110001010010;
    9'd170: Q <= 42'b010010111111000000001000111000011110010000;
    9'd171: Q <= 42'b101011011010010110011101000001111011111001;
    9'd172: Q <= 42'b101010010111001010111011000010110010110100;
    9'd173: Q <= 42'b001000111000110001111010010000010100000010;
    9'd174: Q <= 42'b010011110001111011001000110001001001111010;
    9'd175: Q <= 42'b010000101010110111000111000010010011110001;
    9'd176: Q <= 42'b101010000100110110001000100100011010101010;
    9'd177: Q <= 42'b011000100111101001001110010101101001101011;
    9'd178: Q <= 42'b100101001100001011000011001010000100100100;
    9'd179: Q <= 42'b000010010000110011010110111010111100101001;
    9'd180: Q <= 42'b011000101100110100000111010000100010100101;
    9'd181: Q <= 42'b100010110110010000101010010101010111110010;
    9'd182: Q <= 42'b011111100000110110000101101000110000010010;
    9'd183: Q <= 42'b010000100011100110010000111100110110101110;
    9'd184: Q <= 42'b101101111001011000101111100101110001001110;
    9'd185: Q <= 42'b001101000111110001100010101101110010000110;
    9'd186: Q <= 42'b001110010111101001100011100000110100100000;
    9'd187: Q <= 42'b010100010110011011100101001000111011100000;
    9'd188: Q <= 42'b101000011110010101110001001001010000001111;
    9'd189: Q <= 42'b001100010110110001010010101101100011110101;
    9'd190: Q <= 42'b000101011011011011111100110100010111100010;
    9'd191: Q <= 42'b010111111011111001010011001110110100010010;
    9'd192: Q <= 42'b010001001101000011000110011001011001000111;
    9'd193: Q <= 42'b000111001000100011110111010110111000111111;
    9'd194: Q <= 42'b000100011100000000001001011110111000000011;
    9'd195: Q <= 42'b010001100010011001001110101010110110111111;
    9'd196: Q <= 42'b001110011111001001111011001000101000111110;
    9'd197: Q <= 42'b100000011110101001000010110010010010000000;
    9'd198: Q <= 42'b000101100010010100101010111001001011110111;
    9'd199: Q <= 42'b011001001101100110100010011100010101111110;
    9'd200: Q <= 42'b011110011010000101101111111000110010100000;
    9'd201: Q <= 42'b010011001111001011100101110000111011111101;
    9'd202: Q <= 42'b000101001011110011100001001010110111001010;
    9'd203: Q <= 42'b000011111101101000000001000101000010110001;
    9'd204: Q <= 42'b001111011001100101111011010001011000011110;
    9'd205: Q <= 42'b001110101000000111111000110001010111100100;
    9'd206: Q <= 42'b010011111011100010001111111010001001101001;
    9'd207: Q <= 42'b001001111000000000011111100010000010011001;
    9'd208: Q <= 42'b011010001011011011011010010000010011110001;
    9'd209: Q <= 42'b001010100111011000011111000100001101001100;
    9'd210: Q <= 42'b010110110011000101111011110110110101010111;
    9'd211: Q <= 42'b001100100000000011001011111110000000101111;
    9'd212: Q <= 42'b001000110101000111011111000101111000010011;
    9'd213: Q <= 42'b010001101001100000010010011101010111011110;
    9'd214: Q <= 42'b001010101010100101101000011010101111111100;
    9'd215: Q <= 42'b000100100010000101111101001110000111011001;
    9'd216: Q <= 42'b100111001101000000101000110001011001011100;
    9'd217: Q <= 42'b011011110011110000010100010100110100001111;
    9'd218: Q <= 42'b000000101111011010111000011101001000000000;
    9'd219: Q <= 42'b101100101000001010101000010110011110011010;
    9'd220: Q <= 42'b101001000111101011000100110100000000010100;
    9'd221: Q <= 42'b001001101011101000000101000100100110001010;
    9'd222: Q <= 42'b101001000010101000010100111110011110011101;
    9'd223: Q <= 42'b010000011000100011111110110101001101001011;
    9'd224: Q <= 42'b011110001011001001001001101000111101110111;
    9'd225: Q <= 42'b101010000001110101110110011000101101001110;
    9'd226: Q <= 42'b010110110010001000010111000110011001101010;
    9'd227: Q <= 42'b100000111001000001001000011100010100100010;
    9'd228: Q <= 42'b101001001110111000000011000000111101101011;
    9'd229: Q <= 42'b001011001110011000000001001001001010000011;
    9'd230: Q <= 42'b101011101000010000111001101010111010010101;
    9'd231: Q <= 42'b101100111010101010111101111100010011001010;
    9'd232: Q <= 42'b101111111011000000011011100100101111010100;
    9'd233: Q <= 42'b101011111110110011111100111010101010000000;
    9'd234: Q <= 42'b010010001010011000111011001101000000101010;
    9'd235: Q <= 42'b001110111011010000101100010101010110000101;
    9'd236: Q <= 42'b001011011100010001010010011101000111111101;
    9'd237: Q <= 42'b000011011010100001111010011000110000110001;
    9'd238: Q <= 42'b001001000000110001000101100010010000111000;
    9'd239: Q <= 42'b000000101010100100001110001010010111011001;
    9'd240: Q <= 42'b101101011110010010000001111001010001111110;
    9'd241: Q <= 42'b000110001001010100001001000010001010110010;
    9'd242: Q <= 42'b101110000010110110000101000010010000011111;
    9'd243: Q <= 42'b001110110100011000100000111100010110111100;
    9'd244: Q <= 42'b001010001010101011001011111000100110110011;
    9'd245: Q <= 42'b011011011001100011010000000100000111111010;
    9'd246: Q <= 42'b000111111100111011110101100100100010100100;
    9'd247: Q <= 42'b101011000111100100001100101001011010011000;
    9'd248: Q <= 42'b101000101001110010101000010010001100110101;
    9'd249: Q <= 42'b010010111000100110000001011110100011010101;
    9'd250: Q <= 42'b011111111100000110111100000100000101111001;
    9'd251: Q <= 42'b100100111101011001100000011010111001111001;
    9'd252: Q <= 42'b001111000000001010110101000100000101110111;
    9'd253: Q <= 42'b011101010111110101110100100100101011011000;
    9'd254: Q <= 42'b011001110110001010000101011110001010110001;
    9'd255: Q <= 42'b010100101001110111000000111100110110110111;
    9'd256: Q <= 42'b011010111000110001100011101010010111110010;
    9'd257: Q <= 42'b001101011110110001010101000010101111110011;
    9'd258: Q <= 42'b011001011011000110000001101001100000110101;
    9'd259: Q <= 42'b101011001010000011110111010001100000111100;
    9'd260: Q <= 42'b100101101011100101001011000110010100010001;
    9'd261: Q <= 42'b000111001110010010011001101110111100010010;
    9'd262: Q <= 42'b011111001101000011100100100001010101011000;
    9'd263: Q <= 42'b100011001111010000101010101101000111001010;
    9'd264: Q <= 42'b000001110010011011111100000101110111000011;
    9'd265: Q <= 42'b011110011010011000111100111001110011010000;
    9'd266: Q <= 42'b001101111110101001000001001110011100001110;
    9'd267: Q <= 42'b000010000100101010010010111001111101110110;
    9'd268: Q <= 42'b100010011101110110101001001100110101000001;
    9'd269: Q <= 42'b101100100100101010011110001100000010010010;
    9'd270: Q <= 42'b010000011110101001000111110100011100001100;
    9'd271: Q <= 42'b000011110101100101101001011000000110010110;
    9'd272: Q <= 42'b100010100000111001100011101001100000110011;
    9'd273: Q <= 42'b101000000000110111101011000000001001111100;
    9'd274: Q <= 42'b001100111101010011101111101010100100111000;
    9'd275: Q <= 42'b100100011101000110001110001000101110000011;
    9'd276: Q <= 42'b000000100010110110110111100001100111011001;
    9'd277: Q <= 42'b000000101101000111101000111001101101100110;
    9'd278: Q <= 42'b101010100000000110100110000010100010100111;
    9'd279: Q <= 42'b011110000001000111010100110001101011011111;
    9'd280: Q <= 42'b000000110011000100101000110110100000001110;
    9'd281: Q <= 42'b010010100000110101111110011000110101111011;
    9'd282: Q <= 42'b100100001011010001001010011010010110101110;
    9'd283: Q <= 42'b011010011100111000010001011101000100011010;
    9'd284: Q <= 42'b101110100101011001011000011001011010010101;
    9'd285: Q <= 42'b101010010001010100010110000101100111011000;
    9'd286: Q <= 42'b101010110000011011110110111000001110110000;
    9'd287: Q <= 42'b100010101100100110101011000101110111001000;
    9'd288: Q <= 42'b100110010011101000010011010001101101011010;
    9'd289: Q <= 42'b101011001011010011110001010010010011110101;
    9'd290: Q <= 42'b001100001100010111100100100100000001001000;
    9'd291: Q <= 42'b011011100000110101010100010101110100011111;
    9'd292: Q <= 42'b000100001000011010111110011110000100000001;
    9'd293: Q <= 42'b010101110111100000101000111010101111111011;
    9'd294: Q <= 42'b011001101001010001101010011000101101110001;
    9'd295: Q <= 42'b101000100111010011011110110100011010010001;
    9'd296: Q <= 42'b101011111111000001111100001101110111011000;
    9'd297: Q <= 42'b101010110111110101111111100010101110100001;
    9'd298: Q <= 42'b011001110001110110101101101000101100001011;
    9'd299: Q <= 42'b001011010011100110010001101101100101010001;
    9'd300: Q <= 42'b100000100101101000011100011000001100010111;
    9'd301: Q <= 42'b010111010001110110100110100010111000001011;
    9'd302: Q <= 42'b001001100010100011000111111110000011111011;
    9'd303: Q <= 42'b100000100010100101000101011010100010010100;
    9'd304: Q <= 42'b010011111110111011111100100110000100110000;
    9'd305: Q <= 42'b001101000011110100110101010000000010101010;
    9'd306: Q <= 42'b101111111011010000011001000001000011000001;
    9'd307: Q <= 42'b000101111100100110000000100010110010010111;
    9'd308: Q <= 42'b010010000000001010010100000100001010001000;
    9'd309: Q <= 42'b101110011010110100111101011100100110101110;
    9'd310: Q <= 42'b000101011110110010000111100101111000101100;
    9'd311: Q <= 42'b000000100100101000110100001100101111001011;
    9'd312: Q <= 42'b010111110011101011011111011100011011110111;
    9'd313: Q <= 42'b001101001011111010110000001100000010111101;
    9'd314: Q <= 42'b011100110100000001111011010100101001110000;
    9'd315: Q <= 42'b100010110000001001101101100100100010100001;
    9'd316: Q <= 42'b001110111100010110100011101100001101100001;
    9'd317: Q <= 42'b101111000100100111110001110100010010001000;
    9'd318: Q <= 42'b010010001111101000000001011001010100100011;
    9'd319: Q <= 42'b000011111000100100110011010001111001011011;
    9'd320: Q <= 42'b010101010110000101001100001100100011001101;
    9'd321: Q <= 42'b100100011111101000100100011110000011100100;
    9'd322: Q <= 42'b101101100100110101110010010100010101000110;
    9'd323: Q <= 42'b000010011111001010111111000000010111111010;
    9'd324: Q <= 42'b010110001010001011000000011100011011000110;
    9'd325: Q <= 42'b010001111000100101001101101110110010010010;
    9'd326: Q <= 42'b101000110101010011100111111010001010000011;
    9'd327: Q <= 42'b101110100010100101010100011010011100011101;
    9'd328: Q <= 42'b100111011110000101111100110101111110000111;
    9'd329: Q <= 42'b000001111110101010000001000000110111111010;
    9'd330: Q <= 42'b001100110011000011110010011100001100001010;
    9'd331: Q <= 42'b000101011100001000000110001100011010100101;
    9'd332: Q <= 42'b001000101001000001111000001010110111101111;
    9'd333: Q <= 42'b010111110001010000011101010010001100111101;
    9'd334: Q <= 42'b100111010010100000010011110001111001010110;
    9'd335: Q <= 42'b101011111100111000000110110110100011001000;
    9'd336: Q <= 42'b001010111100001011101000001110111000111000;
    9'd337: Q <= 42'b101000011010111010101011001010010001110100;
    9'd338: Q <= 42'b001010110110000000111100110110011000011101;
    9'd339: Q <= 42'b001010000011110110101100011000011111111110;
    9'd340: Q <= 42'b011010100110111010110001101110111101110110;
    endcase end         
    end
endmodule
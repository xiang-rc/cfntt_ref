module tf_ROM 
    #(parameter addr_rom_width = 10,
                 data_width = 14,
                 depth_rom = 1023)
    (
    input clk,
    input [addr_rom_width-1:0] A,
    input REN,
    output reg [data_width-1:0] Q
    );
    
    always@(posedge clk)
    begin
    if(REN == 1'b1) begin
    case(A)
    10'd0: Q <= 14'd10810;
    10'd1: Q <= 14'd7143;
    10'd2: Q <= 14'd4043;
    10'd3: Q <= 14'd10984;
    10'd4: Q <= 14'd722;
    10'd5: Q <= 14'd5736;
    10'd6: Q <= 14'd8155;
    10'd7: Q <= 14'd3542;
    10'd8: Q <= 14'd8785;
    10'd9: Q <= 14'd9744;
    10'd10: Q <= 14'd3621;
    10'd11: Q <= 14'd10643;
    10'd12: Q <= 14'd1212;
    10'd13: Q <= 14'd3195;
    10'd14: Q <= 14'd5860;
    10'd15: Q <= 14'd7468;
    10'd16: Q <= 14'd2639;
    10'd17: Q <= 14'd9664;
    10'd18: Q <= 14'd11340;
    10'd19: Q <= 14'd11726;
    10'd20: Q <= 14'd9314;
    10'd21: Q <= 14'd9283;
    10'd22: Q <= 14'd9545;
    10'd23: Q <= 14'd5728;
    10'd24: Q <= 14'd7698;
    10'd25: Q <= 14'd5023;
    10'd26: Q <= 14'd5828;
    10'd27: Q <= 14'd8961;
    10'd28: Q <= 14'd6512;
    10'd29: Q <= 14'd7311;
    10'd30: Q <= 14'd1351;
    10'd31: Q <= 14'd2319;
    10'd32: Q <= 14'd11119;
    10'd33: Q <= 14'd11334;
    10'd34: Q <= 14'd11499;
    10'd35: Q <= 14'd9088;
    10'd36: Q <= 14'd3014;
    10'd37: Q <= 14'd5086;
    10'd38: Q <= 14'd10963;
    10'd39: Q <= 14'd4846;
    10'd40: Q <= 14'd9542;
    10'd41: Q <= 14'd9154;
    10'd42: Q <= 14'd3712;
    10'd43: Q <= 14'd4805;
    10'd44: Q <= 14'd8736;
    10'd45: Q <= 14'd11227;
    10'd46: Q <= 14'd9995;
    10'd47: Q <= 14'd3091;
    10'd48: Q <= 14'd12208;
    10'd49: Q <= 14'd7969;
    10'd50: Q <= 14'd11289;
    10'd51: Q <= 14'd9326;
    10'd52: Q <= 14'd7393;
    10'd53: Q <= 14'd9238;
    10'd54: Q <= 14'd2366;
    10'd55: Q <= 14'd11112;
    10'd56: Q <= 14'd8034;
    10'd57: Q <= 14'd10654;
    10'd58: Q <= 14'd9521;
    10'd59: Q <= 14'd12149;
    10'd60: Q <= 14'd10436;
    10'd61: Q <= 14'd7678;
    10'd62: Q <= 14'd11563;
    10'd63: Q <= 14'd1260;
    10'd64: Q <= 14'd4388;
    10'd65: Q <= 14'd4632;
    10'd66: Q <= 14'd6534;
    10'd67: Q <= 14'd2426;
    10'd68: Q <= 14'd334;
    10'd69: Q <= 14'd1428;
    10'd70: Q <= 14'd1696;
    10'd71: Q <= 14'd2013;
    10'd72: Q <= 14'd9000;
    10'd73: Q <= 14'd729;
    10'd74: Q <= 14'd3241;
    10'd75: Q <= 14'd2881;
    10'd76: Q <= 14'd3284;
    10'd77: Q <= 14'd7197;
    10'd78: Q <= 14'd10200;
    10'd79: Q <= 14'd8595;
    10'd80: Q <= 14'd7110;
    10'd81: Q <= 14'd10530;
    10'd82: Q <= 14'd8582;
    10'd83: Q <= 14'd3382;
    10'd84: Q <= 14'd11934;
    10'd85: Q <= 14'd9741;
    10'd86: Q <= 14'd8058;
    10'd87: Q <= 14'd3637;
    10'd88: Q <= 14'd3459;
    10'd89: Q <= 14'd145;
    10'd90: Q <= 14'd6747;
    10'd91: Q <= 14'd9558;
    10'd92: Q <= 14'd8357;
    10'd93: Q <= 14'd7399;
    10'd94: Q <= 14'd6378;
    10'd95: Q <= 14'd9447;
    10'd96: Q <= 14'd480;
    10'd97: Q <= 14'd1022;
    10'd98: Q <= 14'd9;
    10'd99: Q <= 14'd9821;
    10'd100: Q <= 14'd339;
    10'd101: Q <= 14'd5791;
    10'd102: Q <= 14'd544;
    10'd103: Q <= 14'd10616;
    10'd104: Q <= 14'd4278;
    10'd105: Q <= 14'd6958;
    10'd106: Q <= 14'd7300;
    10'd107: Q <= 14'd8112;
    10'd108: Q <= 14'd8705;
    10'd109: Q <= 14'd1381;
    10'd110: Q <= 14'd9764;
    10'd111: Q <= 14'd11336;
    10'd112: Q <= 14'd8541;
    10'd113: Q <= 14'd827;
    10'd114: Q <= 14'd5767;
    10'd115: Q <= 14'd2476;
    10'd116: Q <= 14'd118;
    10'd117: Q <= 14'd2197;
    10'd118: Q <= 14'd7222;
    10'd119: Q <= 14'd3949;
    10'd120: Q <= 14'd8993;
    10'd121: Q <= 14'd4452;
    10'd122: Q <= 14'd2396;
    10'd123: Q <= 14'd7935;
    10'd124: Q <= 14'd130;
    10'd125: Q <= 14'd2837;
    10'd126: Q <= 14'd6915;
    10'd127: Q <= 14'd2401;
    10'd128: Q <= 14'd442;
    10'd129: Q <= 14'd7188;
    10'd130: Q <= 14'd11222;
    10'd131: Q <= 14'd390;
    10'd132: Q <= 14'd773;
    10'd133: Q <= 14'd8456;
    10'd134: Q <= 14'd3778;
    10'd135: Q <= 14'd354;
    10'd136: Q <= 14'd4861;
    10'd137: Q <= 14'd9377;
    10'd138: Q <= 14'd5698;
    10'd139: Q <= 14'd5012;
    10'd140: Q <= 14'd9808;
    10'd141: Q <= 14'd2859;
    10'd142: Q <= 14'd11244;
    10'd143: Q <= 14'd1017;
    10'd144: Q <= 14'd7404;
    10'd145: Q <= 14'd1632;
    10'd146: Q <= 14'd7205;
    10'd147: Q <= 14'd27;
    10'd148: Q <= 14'd9223;
    10'd149: Q <= 14'd8526;
    10'd150: Q <= 14'd10849;
    10'd151: Q <= 14'd1537;
    10'd152: Q <= 14'd242;
    10'd153: Q <= 14'd4714;
    10'd154: Q <= 14'd8146;
    10'd155: Q <= 14'd9611;
    10'd156: Q <= 14'd3704;
    10'd157: Q <= 14'd5019;
    10'd158: Q <= 14'd11744;
    10'd159: Q <= 14'd1002;
    10'd160: Q <= 14'd5011;
    10'd161: Q <= 14'd5088;
    10'd162: Q <= 14'd8005;
    10'd163: Q <= 14'd7313;
    10'd164: Q <= 14'd10682;
    10'd165: Q <= 14'd8509;
    10'd166: Q <= 14'd11414;
    10'd167: Q <= 14'd9852;
    10'd168: Q <= 14'd3646;
    10'd169: Q <= 14'd6022;
    10'd170: Q <= 14'd2987;
    10'd171: Q <= 14'd9723;
    10'd172: Q <= 14'd10102;
    10'd173: Q <= 14'd6250;
    10'd174: Q <= 14'd9867;
    10'd175: Q <= 14'd11224;
    10'd176: Q <= 14'd2143;
    10'd177: Q <= 14'd11885;
    10'd178: Q <= 14'd7644;
    10'd179: Q <= 14'd1168;
    10'd180: Q <= 14'd5277;
    10'd181: Q <= 14'd11082;
    10'd182: Q <= 14'd3248;
    10'd183: Q <= 14'd493;
    10'd184: Q <= 14'd8193;
    10'd185: Q <= 14'd6845;
    10'd186: Q <= 14'd2381;
    10'd187: Q <= 14'd7952;
    10'd188: Q <= 14'd11854;
    10'd189: Q <= 14'd1378;
    10'd190: Q <= 14'd1912;
    10'd191: Q <= 14'd2166;
    10'd192: Q <= 14'd3915;
    10'd193: Q <= 14'd12176;
    10'd194: Q <= 14'd7370;
    10'd195: Q <= 14'd12129;
    10'd196: Q <= 14'd3149;
    10'd197: Q <= 14'd12286;
    10'd198: Q <= 14'd4437;
    10'd199: Q <= 14'd3636;
    10'd200: Q <= 14'd4938;
    10'd201: Q <= 14'd5291;
    10'd202: Q <= 14'd2704;
    10'd203: Q <= 14'd10863;
    10'd204: Q <= 14'd7635;
    10'd205: Q <= 14'd1663;
    10'd206: Q <= 14'd10512;
    10'd207: Q <= 14'd3364;
    10'd208: Q <= 14'd1689;
    10'd209: Q <= 14'd4057;
    10'd210: Q <= 14'd9018;
    10'd211: Q <= 14'd9442;
    10'd212: Q <= 14'd7875;
    10'd213: Q <= 14'd2174;
    10'd214: Q <= 14'd4372;
    10'd215: Q <= 14'd7247;
    10'd216: Q <= 14'd9984;
    10'd217: Q <= 14'd4053;
    10'd218: Q <= 14'd2645;
    10'd219: Q <= 14'd5195;
    10'd220: Q <= 14'd9509;
    10'd221: Q <= 14'd7394;
    10'd222: Q <= 14'd1484;
    10'd223: Q <= 14'd9042;
    10'd224: Q <= 14'd9603;
    10'd225: Q <= 14'd8311;
    10'd226: Q <= 14'd9320;
    10'd227: Q <= 14'd9919;
    10'd228: Q <= 14'd2865;
    10'd229: Q <= 14'd5332;
    10'd230: Q <= 14'd3510;
    10'd231: Q <= 14'd1630;
    10'd232: Q <= 14'd10163;
    10'd233: Q <= 14'd5407;
    10'd234: Q <= 14'd3186;
    10'd235: Q <= 14'd11136;
    10'd236: Q <= 14'd9405;
    10'd237: Q <= 14'd10040;
    10'd238: Q <= 14'd8241;
    10'd239: Q <= 14'd9890;
    10'd240: Q <= 14'd8889;
    10'd241: Q <= 14'd7098;
    10'd242: Q <= 14'd9153;
    10'd243: Q <= 14'd9289;
    10'd244: Q <= 14'd671;
    10'd245: Q <= 14'd3016;
    10'd246: Q <= 14'd243;
    10'd247: Q <= 14'd6730;
    10'd248: Q <= 14'd420;
    10'd249: Q <= 14'd10111;
    10'd250: Q <= 14'd1544;
    10'd251: Q <= 14'd3985;
    10'd252: Q <= 14'd4905;
    10'd253: Q <= 14'd3531;
    10'd254: Q <= 14'd476;
    10'd255: Q <= 14'd49;
    10'd256: Q <= 14'd1263;
    10'd257: Q <= 14'd5915;
    10'd258: Q <= 14'd1483;
    10'd259: Q <= 14'd9789;
    10'd260: Q <= 14'd10800;
    10'd261: Q <= 14'd10706;
    10'd262: Q <= 14'd6347;
    10'd263: Q <= 14'd1512;
    10'd264: Q <= 14'd350;
    10'd265: Q <= 14'd10474;
    10'd266: Q <= 14'd5383;
    10'd267: Q <= 14'd5369;
    10'd268: Q <= 14'd10232;
    10'd269: Q <= 14'd9087;
    10'd270: Q <= 14'd4493;
    10'd271: Q <= 14'd9551;
    10'd272: Q <= 14'd6421;
    10'd273: Q <= 14'd6554;
    10'd274: Q <= 14'd2655;
    10'd275: Q <= 14'd9280;
    10'd276: Q <= 14'd1693;
    10'd277: Q <= 14'd174;
    10'd278: Q <= 14'd723;
    10'd279: Q <= 14'd10314;
    10'd280: Q <= 14'd8532;
    10'd281: Q <= 14'd347;
    10'd282: Q <= 14'd2925;
    10'd283: Q <= 14'd8974;
    10'd284: Q <= 14'd11863;
    10'd285: Q <= 14'd1858;
    10'd286: Q <= 14'd4754;
    10'd287: Q <= 14'd3030;
    10'd288: Q <= 14'd4115;
    10'd289: Q <= 14'd2361;
    10'd290: Q <= 14'd10446;
    10'd291: Q <= 14'd2908;
    10'd292: Q <= 14'd218;
    10'd293: Q <= 14'd3434;
    10'd294: Q <= 14'd8760;
    10'd295: Q <= 14'd3963;
    10'd296: Q <= 14'd576;
    10'd297: Q <= 14'd6142;
    10'd298: Q <= 14'd9842;
    10'd299: Q <= 14'd1954;
    10'd300: Q <= 14'd10238;
    10'd301: Q <= 14'd9407;
    10'd302: Q <= 14'd10484;
    10'd303: Q <= 14'd3991;
    10'd304: Q <= 14'd8320;
    10'd305: Q <= 14'd9522;
    10'd306: Q <= 14'd156;
    10'd307: Q <= 14'd2281;
    10'd308: Q <= 14'd5876;
    10'd309: Q <= 14'd10258;
    10'd310: Q <= 14'd5333;
    10'd311: Q <= 14'd3772;
    10'd312: Q <= 14'd418;
    10'd313: Q <= 14'd5908;
    10'd314: Q <= 14'd11836;
    10'd315: Q <= 14'd5429;
    10'd316: Q <= 14'd7515;
    10'd317: Q <= 14'd7552;
    10'd318: Q <= 14'd1293;
    10'd319: Q <= 14'd295;
    10'd320: Q <= 14'd6099;
    10'd321: Q <= 14'd5766;
    10'd322: Q <= 14'd652;
    10'd323: Q <= 14'd8273;
    10'd324: Q <= 14'd4077;
    10'd325: Q <= 14'd8527;
    10'd326: Q <= 14'd9370;
    10'd327: Q <= 14'd325;
    10'd328: Q <= 14'd10885;
    10'd329: Q <= 14'd11143;
    10'd330: Q <= 14'd11341;
    10'd331: Q <= 14'd5990;
    10'd332: Q <= 14'd1159;
    10'd333: Q <= 14'd8561;
    10'd334: Q <= 14'd8240;
    10'd335: Q <= 14'd3329;
    10'd336: Q <= 14'd4298;
    10'd337: Q <= 14'd12121;
    10'd338: Q <= 14'd2692;
    10'd339: Q <= 14'd5961;
    10'd340: Q <= 14'd7183;
    10'd341: Q <= 14'd10327;
    10'd342: Q <= 14'd1594;
    10'd343: Q <= 14'd6167;
    10'd344: Q <= 14'd9734;
    10'd345: Q <= 14'd7105;
    10'd346: Q <= 14'd11089;
    10'd347: Q <= 14'd1360;
    10'd348: Q <= 14'd3956;
    10'd349: Q <= 14'd6170;
    10'd350: Q <= 14'd5297;
    10'd351: Q <= 14'd8210;
    10'd352: Q <= 14'd11231;
    10'd353: Q <= 14'd922;
    10'd354: Q <= 14'd441;
    10'd355: Q <= 14'd1958;
    10'd356: Q <= 14'd4322;
    10'd357: Q <= 14'd1112;
    10'd358: Q <= 14'd2078;
    10'd359: Q <= 14'd4046;
    10'd360: Q <= 14'd709;
    10'd361: Q <= 14'd9139;
    10'd362: Q <= 14'd1319;
    10'd363: Q <= 14'd4240;
    10'd364: Q <= 14'd8719;
    10'd365: Q <= 14'd6224;
    10'd366: Q <= 14'd11454;
    10'd367: Q <= 14'd2459;
    10'd368: Q <= 14'd683;
    10'd369: Q <= 14'd3656;
    10'd370: Q <= 14'd12225;
    10'd371: Q <= 14'd10723;
    10'd372: Q <= 14'd5782;
    10'd373: Q <= 14'd9341;
    10'd374: Q <= 14'd9786;
    10'd375: Q <= 14'd9166;
    10'd376: Q <= 14'd10542;
    10'd377: Q <= 14'd9235;
    10'd378: Q <= 14'd6803;
    10'd379: Q <= 14'd7856;
    10'd380: Q <= 14'd6370;
    10'd381: Q <= 14'd3834;
    10'd382: Q <= 14'd7032;
    10'd383: Q <= 14'd7048;
    10'd384: Q <= 14'd9369;
    10'd385: Q <= 14'd8120;
    10'd386: Q <= 14'd9162;
    10'd387: Q <= 14'd6821;
    10'd388: Q <= 14'd1010;
    10'd389: Q <= 14'd8807;
    10'd390: Q <= 14'd787;
    10'd391: Q <= 14'd5057;
    10'd392: Q <= 14'd4698;
    10'd393: Q <= 14'd4780;
    10'd394: Q <= 14'd8844;
    10'd395: Q <= 14'd12097;
    10'd396: Q <= 14'd1321;
    10'd397: Q <= 14'd4912;
    10'd398: Q <= 14'd10240;
    10'd399: Q <= 14'd677;
    10'd400: Q <= 14'd6415;
    10'd401: Q <= 14'd6234;
    10'd402: Q <= 14'd8953;
    10'd403: Q <= 14'd1323;
    10'd404: Q <= 14'd9523;
    10'd405: Q <= 14'd12237;
    10'd406: Q <= 14'd3174;
    10'd407: Q <= 14'd1579;
    10'd408: Q <= 14'd11858;
    10'd409: Q <= 14'd9784;
    10'd410: Q <= 14'd5906;
    10'd411: Q <= 14'd3957;
    10'd412: Q <= 14'd9450;
    10'd413: Q <= 14'd151;
    10'd414: Q <= 14'd10162;
    10'd415: Q <= 14'd12231;
    10'd416: Q <= 14'd12048;
    10'd417: Q <= 14'd3532;
    10'd418: Q <= 14'd11286;
    10'd419: Q <= 14'd1956;
    10'd420: Q <= 14'd7280;
    10'd421: Q <= 14'd11404;
    10'd422: Q <= 14'd6281;
    10'd423: Q <= 14'd3477;
    10'd424: Q <= 14'd6608;
    10'd425: Q <= 14'd142;
    10'd426: Q <= 14'd11184;
    10'd427: Q <= 14'd9445;
    10'd428: Q <= 14'd3438;
    10'd429: Q <= 14'd11314;
    10'd430: Q <= 14'd4212;
    10'd431: Q <= 14'd9260;
    10'd432: Q <= 14'd6695;
    10'd433: Q <= 14'd4782;
    10'd434: Q <= 14'd5886;
    10'd435: Q <= 14'd8076;
    10'd436: Q <= 14'd504;
    10'd437: Q <= 14'd2302;
    10'd438: Q <= 14'd11684;
    10'd439: Q <= 14'd11868;
    10'd440: Q <= 14'd8209;
    10'd441: Q <= 14'd3602;
    10'd442: Q <= 14'd6068;
    10'd443: Q <= 14'd8689;
    10'd444: Q <= 14'd3263;
    10'd445: Q <= 14'd6077;
    10'd446: Q <= 14'd7665;
    10'd447: Q <= 14'd7822;
    10'd448: Q <= 14'd7500;
    10'd449: Q <= 14'd6752;
    10'd450: Q <= 14'd4749;
    10'd451: Q <= 14'd4449;
    10'd452: Q <= 14'd6833;
    10'd453: Q <= 14'd12142;
    10'd454: Q <= 14'd8500;
    10'd455: Q <= 14'd6118;
    10'd456: Q <= 14'd8471;
    10'd457: Q <= 14'd1190;
    10'd458: Q <= 14'd9606;
    10'd459: Q <= 14'd3860;
    10'd460: Q <= 14'd5445;
    10'd461: Q <= 14'd7753;
    10'd462: Q <= 14'd11239;
    10'd463: Q <= 14'd5079;
    10'd464: Q <= 14'd9027;
    10'd465: Q <= 14'd2169;
    10'd466: Q <= 14'd11767;
    10'd467: Q <= 14'd7965;
    10'd468: Q <= 14'd4916;
    10'd469: Q <= 14'd8214;
    10'd470: Q <= 14'd5315;
    10'd471: Q <= 14'd11011;
    10'd472: Q <= 14'd9945;
    10'd473: Q <= 14'd1973;
    10'd474: Q <= 14'd6715;
    10'd475: Q <= 14'd8775;
    10'd476: Q <= 14'd11248;
    10'd477: Q <= 14'd5925;
    10'd478: Q <= 14'd11271;
    10'd479: Q <= 14'd654;
    10'd480: Q <= 14'd3565;
    10'd481: Q <= 14'd1702;
    10'd482: Q <= 14'd1987;
    10'd483: Q <= 14'd6760;
    10'd484: Q <= 14'd5206;
    10'd485: Q <= 14'd3199;
    10'd486: Q <= 14'd12233;
    10'd487: Q <= 14'd6136;
    10'd488: Q <= 14'd6427;
    10'd489: Q <= 14'd6874;
    10'd490: Q <= 14'd8646;
    10'd491: Q <= 14'd4948;
    10'd492: Q <= 14'd6152;
    10'd493: Q <= 14'd400;
    10'd494: Q <= 14'd10561;
    10'd495: Q <= 14'd5339;
    10'd496: Q <= 14'd5446;
    10'd497: Q <= 14'd3710;
    10'd498: Q <= 14'd6093;
    10'd499: Q <= 14'd468;
    10'd500: Q <= 14'd8301;
    10'd501: Q <= 14'd316;
    10'd502: Q <= 14'd11907;
    10'd503: Q <= 14'd10256;
    10'd504: Q <= 14'd8291;
    10'd505: Q <= 14'd3879;
    10'd506: Q <= 14'd1922;
    10'd507: Q <= 14'd10930;
    10'd508: Q <= 14'd6854;
    10'd509: Q <= 14'd973;
    10'd510: Q <= 14'd11035;
    10'd511: Q <= 14'd7;
    10'd512: Q <= 14'd1936;
    10'd513: Q <= 14'd845;
    10'd514: Q <= 14'd3723;
    10'd515: Q <= 14'd3154;
    10'd516: Q <= 14'd5054;
    10'd517: Q <= 14'd3285;
    10'd518: Q <= 14'd7929;
    10'd519: Q <= 14'd216;
    10'd520: Q <= 14'd50;
    10'd521: Q <= 14'd6763;
    10'd522: Q <= 14'd769;
    10'd523: Q <= 14'd767;
    10'd524: Q <= 14'd8484;
    10'd525: Q <= 14'd10076;
    10'd526: Q <= 14'd4153;
    10'd527: Q <= 14'd3120;
    10'd528: Q <= 14'd6184;
    10'd529: Q <= 14'd6203;
    10'd530: Q <= 14'd5646;
    10'd531: Q <= 14'd8348;
    10'd532: Q <= 14'd3753;
    10'd533: Q <= 14'd3536;
    10'd534: Q <= 14'd5370;
    10'd535: Q <= 14'd3229;
    10'd536: Q <= 14'd4730;
    10'd537: Q <= 14'd10583;
    10'd538: Q <= 14'd3929;
    10'd539: Q <= 14'd1282;
    10'd540: Q <= 14'd8717;
    10'd541: Q <= 14'd2021;
    10'd542: Q <= 14'd9457;
    10'd543: Q <= 14'd3944;
    10'd544: Q <= 14'd4099;
    10'd545: Q <= 14'd5604;
    10'd546: Q <= 14'd6759;
    10'd547: Q <= 14'd2171;
    10'd548: Q <= 14'd8809;
    10'd549: Q <= 14'd11024;
    10'd550: Q <= 14'd3007;
    10'd551: Q <= 14'd9344;
    10'd552: Q <= 14'd5349;
    10'd553: Q <= 14'd2633;
    10'd554: Q <= 14'd1406;
    10'd555: Q <= 14'd9057;
    10'd556: Q <= 14'd11996;
    10'd557: Q <= 14'd4855;
    10'd558: Q <= 14'd8520;
    10'd559: Q <= 14'd9348;
    10'd560: Q <= 14'd11722;
    10'd561: Q <= 14'd6627;
    10'd562: Q <= 14'd5289;
    10'd563: Q <= 14'd3837;
    10'd564: Q <= 14'd2595;
    10'd565: Q <= 14'd3221;
    10'd566: Q <= 14'd4273;
    10'd567: Q <= 14'd4050;
    10'd568: Q <= 14'd7082;
    10'd569: Q <= 14'd844;
    10'd570: Q <= 14'd5202;
    10'd571: Q <= 14'd11309;
    10'd572: Q <= 14'd11607;
    10'd573: Q <= 14'd4590;
    10'd574: Q <= 14'd7207;
    10'd575: Q <= 14'd8820;
    10'd576: Q <= 14'd6138;
    10'd577: Q <= 14'd7846;
    10'd578: Q <= 14'd8871;
    10'd579: Q <= 14'd4693;
    10'd580: Q <= 14'd2338;
    10'd581: Q <= 14'd9996;
    10'd582: Q <= 14'd11872;
    10'd583: Q <= 14'd1802;
    10'd584: Q <= 14'd1555;
    10'd585: Q <= 14'd5103;
    10'd586: Q <= 14'd10398;
    10'd587: Q <= 14'd7878;
    10'd588: Q <= 14'd10699;
    10'd589: Q <= 14'd1223;
    10'd590: Q <= 14'd9955;
    10'd591: Q <= 14'd11009;
    10'd592: Q <= 14'd614;
    10'd593: Q <= 14'd12265;
    10'd594: Q <= 14'd10918;
    10'd595: Q <= 14'd11385;
    10'd596: Q <= 14'd9804;
    10'd597: Q <= 14'd6742;
    10'd598: Q <= 14'd7250;
    10'd599: Q <= 14'd881;
    10'd600: Q <= 14'd11924;
    10'd601: Q <= 14'd1015;
    10'd602: Q <= 14'd10362;
    10'd603: Q <= 14'd5461;
    10'd604: Q <= 14'd9343;
    10'd605: Q <= 14'd2637;
    10'd606: Q <= 14'd7779;
    10'd607: Q <= 14'd4684;
    10'd608: Q <= 14'd3360;
    10'd609: Q <= 14'd7154;
    10'd610: Q <= 14'd63;
    10'd611: Q <= 14'd7302;
    10'd612: Q <= 14'd2373;
    10'd613: Q <= 14'd3670;
    10'd614: Q <= 14'd3808;
    10'd615: Q <= 14'd578;
    10'd616: Q <= 14'd5368;
    10'd617: Q <= 14'd11839;
    10'd618: Q <= 14'd1944;
    10'd619: Q <= 14'd7628;
    10'd620: Q <= 14'd11779;
    10'd621: Q <= 14'd9667;
    10'd622: Q <= 14'd6903;
    10'd623: Q <= 14'd5618;
    10'd624: Q <= 14'd10631;
    10'd625: Q <= 14'd5789;
    10'd626: Q <= 14'd3502;
    10'd627: Q <= 14'd5043;
    10'd628: Q <= 14'd826;
    10'd629: Q <= 14'd3090;
    10'd630: Q <= 14'd1398;
    10'd631: Q <= 14'd3065;
    10'd632: Q <= 14'd1506;
    10'd633: Q <= 14'd6586;
    10'd634: Q <= 14'd4483;
    10'd635: Q <= 14'd6389;
    10'd636: Q <= 14'd910;
    10'd637: Q <= 14'd7570;
    10'd638: Q <= 14'd11538;
    10'd639: Q <= 14'd4518;
    10'd640: Q <= 14'd3094;
    10'd641: Q <= 14'd1160;
    10'd642: Q <= 14'd4820;
    10'd643: Q <= 14'd2730;
    10'd644: Q <= 14'd5411;
    10'd645: Q <= 14'd10036;
    10'd646: Q <= 14'd1868;
    10'd647: Q <= 14'd2478;
    10'd648: Q <= 14'd9449;
    10'd649: Q <= 14'd4194;
    10'd650: Q <= 14'd3019;
    10'd651: Q <= 14'd10506;
    10'd652: Q <= 14'd7211;
    10'd653: Q <= 14'd7724;
    10'd654: Q <= 14'd4974;
    10'd655: Q <= 14'd7119;
    10'd656: Q <= 14'd2672;
    10'd657: Q <= 14'd11424;
    10'd658: Q <= 14'd1279;
    10'd659: Q <= 14'd189;
    10'd660: Q <= 14'd3116;
    10'd661: Q <= 14'd10526;
    10'd662: Q <= 14'd2209;
    10'd663: Q <= 14'd10759;
    10'd664: Q <= 14'd1694;
    10'd665: Q <= 14'd8420;
    10'd666: Q <= 14'd7866;
    10'd667: Q <= 14'd5832;
    10'd668: Q <= 14'd1350;
    10'd669: Q <= 14'd10555;
    10'd670: Q <= 14'd8474;
    10'd671: Q <= 14'd7014;
    10'd672: Q <= 14'd10499;
    10'd673: Q <= 14'd11038;
    10'd674: Q <= 14'd6879;
    10'd675: Q <= 14'd2035;
    10'd676: Q <= 14'd1040;
    10'd677: Q <= 14'd10407;
    10'd678: Q <= 14'd6164;
    10'd679: Q <= 14'd7519;
    10'd680: Q <= 14'd944;
    10'd681: Q <= 14'd5287;
    10'd682: Q <= 14'd8620;
    10'd683: Q <= 14'd6616;
    10'd684: Q <= 14'd9269;
    10'd685: Q <= 14'd6883;
    10'd686: Q <= 14'd7624;
    10'd687: Q <= 14'd4834;
    10'd688: Q <= 14'd2712;
    10'd689: Q <= 14'd9461;
    10'd690: Q <= 14'd4352;
    10'd691: Q <= 14'd8176;
    10'd692: Q <= 14'd72;
    10'd693: Q <= 14'd3840;
    10'd694: Q <= 14'd10447;
    10'd695: Q <= 14'd3451;
    10'd696: Q <= 14'd8195;
    10'd697: Q <= 14'd11048;
    10'd698: Q <= 14'd4378;
    10'd699: Q <= 14'd6508;
    10'd700: Q <= 14'd9244;
    10'd701: Q <= 14'd9646;
    10'd702: Q <= 14'd1095;
    10'd703: Q <= 14'd2873;
    10'd704: Q <= 14'd2827;
    10'd705: Q <= 14'd11498;
    10'd706: Q <= 14'd2434;
    10'd707: Q <= 14'd11169;
    10'd708: Q <= 14'd9754;
    10'd709: Q <= 14'd12268;
    10'd710: Q <= 14'd6481;
    10'd711: Q <= 14'd874;
    10'd712: Q <= 14'd9988;
    10'd713: Q <= 14'd170;
    10'd714: Q <= 14'd6639;
    10'd715: Q <= 14'd2307;
    10'd716: Q <= 14'd4289;
    10'd717: Q <= 14'd11641;
    10'd718: Q <= 14'd12139;
    10'd719: Q <= 14'd11259;
    10'd720: Q <= 14'd11823;
    10'd721: Q <= 14'd3821;
    10'd722: Q <= 14'd1681;
    10'd723: Q <= 14'd4649;
    10'd724: Q <= 14'd5969;
    10'd725: Q <= 14'd2929;
    10'd726: Q <= 14'd6026;
    10'd727: Q <= 14'd1573;
    10'd728: Q <= 14'd8443;
    10'd729: Q <= 14'd3793;
    10'd730: Q <= 14'd6226;
    10'd731: Q <= 14'd11787;
    10'd732: Q <= 14'd5118;
    10'd733: Q <= 14'd2602;
    10'd734: Q <= 14'd10388;
    10'd735: Q <= 14'd1849;
    10'd736: Q <= 14'd5776;
    10'd737: Q <= 14'd9021;
    10'd738: Q <= 14'd3795;
    10'd739: Q <= 14'd7988;
    10'd740: Q <= 14'd7766;
    10'd741: Q <= 14'd457;
    10'd742: Q <= 14'd12281;
    10'd743: Q <= 14'd11410;
    10'd744: Q <= 14'd9696;
    10'd745: Q <= 14'd982;
    10'd746: Q <= 14'd10013;
    10'd747: Q <= 14'd4218;
    10'd748: Q <= 14'd4390;
    10'd749: Q <= 14'd8835;
    10'd750: Q <= 14'd8531;
    10'd751: Q <= 14'd7785;
    10'd752: Q <= 14'd778;
    10'd753: Q <= 14'd530;
    10'd754: Q <= 14'd2626;
    10'd755: Q <= 14'd3578;
    10'd756: Q <= 14'd4697;
    10'd757: Q <= 14'd8823;
    10'd758: Q <= 14'd1701;
    10'd759: Q <= 14'd10243;
    10'd760: Q <= 14'd2940;
    10'd761: Q <= 14'd9332;
    10'd762: Q <= 14'd10808;
    10'd763: Q <= 14'd3317;
    10'd764: Q <= 14'd9757;
    10'd765: Q <= 14'd139;
    10'd766: Q <= 14'd3332;
    10'd767: Q <= 14'd343;
    10'd768: Q <= 14'd8841;
    10'd769: Q <= 14'd4538;
    10'd770: Q <= 14'd10381;
    10'd771: Q <= 14'd7078;
    10'd772: Q <= 14'd1866;
    10'd773: Q <= 14'd1208;
    10'd774: Q <= 14'd7562;
    10'd775: Q <= 14'd10584;
    10'd776: Q <= 14'd2450;
    10'd777: Q <= 14'd11873;
    10'd778: Q <= 14'd814;
    10'd779: Q <= 14'd716;
    10'd780: Q <= 14'd10179;
    10'd781: Q <= 14'd2164;
    10'd782: Q <= 14'd6873;
    10'd783: Q <= 14'd5412;
    10'd784: Q <= 14'd8080;
    10'd785: Q <= 14'd9011;
    10'd786: Q <= 14'd6296;
    10'd787: Q <= 14'd3515;
    10'd788: Q <= 14'd11851;
    10'd789: Q <= 14'd1218;
    10'd790: Q <= 14'd5061;
    10'd791: Q <= 14'd10753;
    10'd792: Q <= 14'd10568;
    10'd793: Q <= 14'd2429;
    10'd794: Q <= 14'd8186;
    10'd795: Q <= 14'd1373;
    10'd796: Q <= 14'd9307;
    10'd797: Q <= 14'd717;
    10'd798: Q <= 14'd8700;
    10'd799: Q <= 14'd8921;
    10'd800: Q <= 14'd4227;
    10'd801: Q <= 14'd4238;
    10'd802: Q <= 14'd11677;
    10'd803: Q <= 14'd8067;
    10'd804: Q <= 14'd1526;
    10'd805: Q <= 14'd11749;
    10'd806: Q <= 14'd12164;
    10'd807: Q <= 14'd3163;
    10'd808: Q <= 14'd4032;
    10'd809: Q <= 14'd6127;
    10'd810: Q <= 14'd7449;
    10'd811: Q <= 14'd1389;
    10'd812: Q <= 14'd10221;
    10'd813: Q <= 14'd4404;
    10'd814: Q <= 14'd11943;
    10'd815: Q <= 14'd3359;
    10'd816: Q <= 14'd9084;
    10'd817: Q <= 14'd5209;
    10'd818: Q <= 14'd1092;
    10'd819: Q <= 14'd3678;
    10'd820: Q <= 14'd4265;
    10'd821: Q <= 14'd10361;
    10'd822: Q <= 14'd464;
    10'd823: Q <= 14'd1826;
    10'd824: Q <= 14'd2926;
    10'd825: Q <= 14'd4489;
    10'd826: Q <= 14'd9118;
    10'd827: Q <= 14'd1136;
    10'd828: Q <= 14'd3449;
    10'd829: Q <= 14'd3708;
    10'd830: Q <= 14'd9051;
    10'd831: Q <= 14'd2065;
    10'd832: Q <= 14'd5826;
    10'd833: Q <= 14'd3495;
    10'd834: Q <= 14'd4564;
    10'd835: Q <= 14'd8755;
    10'd836: Q <= 14'd3961;
    10'd837: Q <= 14'd10533;
    10'd838: Q <= 14'd4145;
    10'd839: Q <= 14'd2275;
    10'd840: Q <= 14'd2461;
    10'd841: Q <= 14'd4267;
    10'd842: Q <= 14'd5653;
    10'd843: Q <= 14'd5063;
    10'd844: Q <= 14'd8113;
    10'd845: Q <= 14'd10771;
    10'd846: Q <= 14'd8524;
    10'd847: Q <= 14'd11014;
    10'd848: Q <= 14'd5508;
    10'd849: Q <= 14'd11113;
    10'd850: Q <= 14'd6555;
    10'd851: Q <= 14'd4860;
    10'd852: Q <= 14'd1125;
    10'd853: Q <= 14'd10844;
    10'd854: Q <= 14'd11158;
    10'd855: Q <= 14'd6302;
    10'd856: Q <= 14'd6693;
    10'd857: Q <= 14'd579;
    10'd858: Q <= 14'd3889;
    10'd859: Q <= 14'd9520;
    10'd860: Q <= 14'd3114;
    10'd861: Q <= 14'd6323;
    10'd862: Q <= 14'd212;
    10'd863: Q <= 14'd8314;
    10'd864: Q <= 14'd4883;
    10'd865: Q <= 14'd6454;
    10'd866: Q <= 14'd3087;
    10'd867: Q <= 14'd1417;
    10'd868: Q <= 14'd5676;
    10'd869: Q <= 14'd7784;
    10'd870: Q <= 14'd2257;
    10'd871: Q <= 14'd3744;
    10'd872: Q <= 14'd4963;
    10'd873: Q <= 14'd2528;
    10'd874: Q <= 14'd9233;
    10'd875: Q <= 14'd5102;
    10'd876: Q <= 14'd11877;
    10'd877: Q <= 14'd6701;
    10'd878: Q <= 14'd6444;
    10'd879: Q <= 14'd4924;
    10'd880: Q <= 14'd4781;
    10'd881: Q <= 14'd1014;
    10'd882: Q <= 14'd11841;
    10'd883: Q <= 14'd1327;
    10'd884: Q <= 14'd3607;
    10'd885: Q <= 14'd3942;
    10'd886: Q <= 14'd7057;
    10'd887: Q <= 14'd2717;
    10'd888: Q <= 14'd60;
    10'd889: Q <= 14'd3200;
    10'd890: Q <= 14'd10754;
    10'd891: Q <= 14'd5836;
    10'd892: Q <= 14'd7723;
    10'd893: Q <= 14'd2260;
    10'd894: Q <= 14'd68;
    10'd895: Q <= 14'd180;
    10'd896: Q <= 14'd4138;
    10'd897: Q <= 14'd7684;
    10'd898: Q <= 14'd2689;
    10'd899: Q <= 14'd10880;
    10'd900: Q <= 14'd7070;
    10'd901: Q <= 14'd204;
    10'd902: Q <= 14'd5509;
    10'd903: Q <= 14'd10821;
    10'd904: Q <= 14'd8308;
    10'd905: Q <= 14'd8882;
    10'd906: Q <= 14'd463;
    10'd907: Q <= 14'd10945;
    10'd908: Q <= 14'd9247;
    10'd909: Q <= 14'd9806;
    10'd910: Q <= 14'd10235;
    10'd911: Q <= 14'd4739;
    10'd912: Q <= 14'd8038;
    10'd913: Q <= 14'd6771;
    10'd914: Q <= 14'd1226;
    10'd915: Q <= 14'd9261;
    10'd916: Q <= 14'd5216;
    10'd917: Q <= 14'd11925;
    10'd918: Q <= 14'd9929;
    10'd919: Q <= 14'd11053;
    10'd920: Q <= 14'd9272;
    10'd921: Q <= 14'd7043;
    10'd922: Q <= 14'd4475;
    10'd923: Q <= 14'd3121;
    10'd924: Q <= 14'd4705;
    10'd925: Q <= 14'd1057;
    10'd926: Q <= 14'd9689;
    10'd927: Q <= 14'd11883;
    10'd928: Q <= 14'd10602;
    10'd929: Q <= 14'd146;
    10'd930: Q <= 14'd5268;
    10'd931: Q <= 14'd1403;
    10'd932: Q <= 14'd1804;
    10'd933: Q <= 14'd6094;
    10'd934: Q <= 14'd7100;
    10'd935: Q <= 14'd12050;
    10'd936: Q <= 14'd9389;
    10'd937: Q <= 14'd994;
    10'd938: Q <= 14'd4554;
    10'd939: Q <= 14'd4670;
    10'd940: Q <= 14'd11777;
    10'd941: Q <= 14'd5464;
    10'd942: Q <= 14'd4906;
    10'd943: Q <= 14'd3375;
    10'd944: Q <= 14'd9998;
    10'd945: Q <= 14'd8896;
    10'd946: Q <= 14'd4335;
    10'd947: Q <= 14'd7376;
    10'd948: Q <= 14'd3528;
    10'd949: Q <= 14'd3825;
    10'd950: Q <= 14'd8054;
    10'd951: Q <= 14'd9342;
    10'd952: Q <= 14'd8307;
    10'd953: Q <= 14'd636;
    10'd954: Q <= 14'd5609;
    10'd955: Q <= 14'd11667;
    10'd956: Q <= 14'd10552;
    10'd957: Q <= 14'd5672;
    10'd958: Q <= 14'd4499;
    10'd959: Q <= 14'd5598;
    10'd960: Q <= 14'd3344;
    10'd961: Q <= 14'd10397;
    10'd962: Q <= 14'd8665;
    10'd963: Q <= 14'd6565;
    10'd964: Q <= 14'd10964;
    10'd965: Q <= 14'd11260;
    10'd966: Q <= 14'd10344;
    10'd967: Q <= 14'd5959;
    10'd968: Q <= 14'd10141;
    10'd969: Q <= 14'd8330;
    10'd970: Q <= 14'd5797;
    10'd971: Q <= 14'd2442;
    10'd972: Q <= 14'd1248;
    10'd973: Q <= 14'd5115;
    10'd974: Q <= 14'd4939;
    10'd975: Q <= 14'd10975;
    10'd976: Q <= 14'd1744;
    10'd977: Q <= 14'd2894;
    10'd978: Q <= 14'd8635;
    10'd979: Q <= 14'd6599;
    10'd980: Q <= 14'd9834;
    10'd981: Q <= 14'd8342;
    10'd982: Q <= 14'd338;
    10'd983: Q <= 14'd3343;
    10'd984: Q <= 14'd8170;
    10'd985: Q <= 14'd1522;
    10'd986: Q <= 14'd10138;
    10'd987: Q <= 14'd12269;
    10'd988: Q <= 14'd5002;
    10'd989: Q <= 14'd4608;
    10'd990: Q <= 14'd5163;
    10'd991: Q <= 14'd4578;
    10'd992: Q <= 14'd377;
    10'd993: Q <= 14'd11914;
    10'd994: Q <= 14'd1620;
    10'd995: Q <= 14'd10453;
    10'd996: Q <= 14'd11864;
    10'd997: Q <= 14'd10104;
    10'd998: Q <= 14'd11897;
    10'd999: Q <= 14'd6085;
    10'd1000: Q <= 14'd8122;
    10'd1001: Q <= 14'd11251;
    10'd1002: Q <= 14'd11366;
    10'd1003: Q <= 14'd10058;
    10'd1004: Q <= 14'd6197;
    10'd1005: Q <= 14'd2800;
    10'd1006: Q <= 14'd193;
    10'd1007: Q <= 14'd506;
    10'd1008: Q <= 14'd1255;
    10'd1009: Q <= 14'd1392;
    10'd1010: Q <= 14'd5784;
    10'd1011: Q <= 14'd3276;
    10'd1012: Q <= 14'd8951;
    10'd1013: Q <= 14'd2212;
    10'd1014: Q <= 14'd9615;
    10'd1015: Q <= 14'd10347;
    10'd1016: Q <= 14'd8881;
    10'd1017: Q <= 14'd2575;
    10'd1018: Q <= 14'd1165;
    10'd1019: Q <= 14'd2776;
    10'd1020: Q <= 14'd11111;
    10'd1021: Q <= 14'd6811;
    10'd1022: Q <= 14'd3511;
    endcase end         
    end
endmodule